library ieee;
use ieee.std_logic_1164.all;

entity loop0 is port(
  clk    	: in std_logic;
  input   	: in std_logic_vector (7 downto 0);
  dataValid	: in std_logic;
  rst		: in std_logic;
  output	: out std_logic_vector (7 downto 0);
  start		: out std_logic);
end loop0;

architecture behav of loop0 is

begin
clocked : process(clk, rst)
begin
  if (rst = '1') then
    start <= '0';
  elsif (clk'event and clk = '1') then
    if (dataValid = '1') then
      output <= input;
      start <= '1';
    end if;
    start <= '0';
  end if;
end process clocked;
end behav;